library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PC is
    port(
        clk     : in  std_logic;
        reset_n : in  std_logic;
        en      : in  std_logic;
        sel_a   : in  std_logic;
        sel_imm : in  std_logic;
        add_imm : in  std_logic;
        imm     : in  std_logic_vector(15 downto 0);
        a       : in  std_logic_vector(15 downto 0);
        addr    : out std_logic_vector(31 downto 0)
    );
end PC;

architecture synth of PC is

signal s_curr_addr : std_logic_vector(31 downto 0):=X"00000000";
begin

PC_process: process(clk, reset_n)
begin
	if (reset_n ='0') then
		s_curr_addr <= (31 downto 0 => '0');
	elsif rising_edge(clk) then
		if (en='1') then

			--s_curr_addr <= std_logic_vector(unsigned(s_curr_addr) + 4); --ADDED

			-- BRANCH
			if (add_imm = '1') then
			s_curr_addr <= std_logic_vector(signed(s_curr_addr) + signed(imm(15 downto 2) & "00"));
			
			-- CALL & JMPI
			elsif (sel_imm = '1') then
			s_curr_addr <= std_logic_vector(unsigned(X"0000" & imm(13 downto 0) & "00"));

			-- CALLR
			elsif(sel_a='1') then
			s_curr_addr <= std_logic_vector(unsigned(X"0000" & a(15 downto 2) & "00"));
			
			-- ELSE
			else
			s_curr_addr <= std_logic_vector(signed(s_curr_addr) +4 );
			end if; 
			
		end if;
		
	end if;
end process;

addr <= (X"0000" & s_curr_addr(15 downto 0));
end synth;
