library ieee;
use ieee.std_logic_1164.all;

entity ROM is
    port(
        clk     : in  std_logic;
        cs      : in  std_logic;
        read    : in  std_logic;
        address : in  std_logic_vector(9 downto 0);
        rddata  : out std_logic_vector(31 downto 0)
    );
end ROM;

architecture synth of ROM is

COMPONENT ROM_block
	PORT(
		address		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		clock		: IN STD_LOGIC;
		q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT;

signal s_q : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN

rom_Blck : ROM_block
PORT MAP(clock => clk,
		 address => address,
		  q => s_q);



read_process: process(clk)
begin 
	rddata <= (others => 'Z');
	if(rising_edge(clk)) then
		if(cs = '1' and read = '1') then
			rddata <= s_q;
		end if;
		
	end if;
end process;

end synth;
